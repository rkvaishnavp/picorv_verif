class picorv_base_test extends uvm_test;

  picorv_env env;
  `uvm_component_utils(picorv_base_test)
  `new_comp


endclass  //picorv_base_test extends uvm_test
