class pico_base_test extends uvm_test;

  pico_env env;

endclass //pico_base_test extends uvm_test