`ifndef TB_INCLUDES_SVH
`define TB_INCLUDES_SVH

`endif
