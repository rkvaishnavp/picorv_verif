class picorv_base_seq extends uvm_sequence;

  `uvm_object_utils(picorv_base_seq)
  `new_obj
endclass  //picorv_base_seq extends uvm_sequence
