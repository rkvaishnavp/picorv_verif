class pico_env extends uvm_env;



  function new();
    
  endfunction //new()
endclass //pico_env extends uvm_env