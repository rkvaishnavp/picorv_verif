package axil_pkg;
  parameter int DATA_WIDTH = 32;
  parameter int ADDR_WIDTH = 16;
  parameter bit PIPELINE_OUTPUT = 0;
endpackage
