class pico_agent extends uvm_agent;

  

  `uvm_component_utils(pico_agent)
  `new_comp

endclass //pico_agent extends uvm_agent